`define DATA_WIDTH 8
`define CMD_WIDTH 4

`define num_transaction 10

`define SHIFT_WIDTH  $clog2(`DATA_WIDTH)
