`define DATA_WIDTH 16
`define CMD_WIDTH 4

`define num_transactions 20

parameter POW_2_N = $clog2(`DATA_WIDTH);
