`define DATA_WIDTH 16
`define CMD_WIDTH 4

`define num_transactions 20
